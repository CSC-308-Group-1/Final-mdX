//////////////////////////////////////////////////////////////////////////////////////////
//    ENGR_850 Term Project
//    File        : Defines.sv
//    Authors     : Arok Lijo J , Chandan Gireesha , Saifulla 
//    Description : Testbench Defines
//////////////////////////////////////////////////////////////////////////////////////////

`define SMEM_MAX 1024
`define RMEM_MAX 256
`define TRANSACTION_COUNT 800
`define DRIV_IF mem_intf.ME_DRIVER.ME_driver_cb
`define MON_IF mem_intf.ME_MONITOR.ME_monitor_cb