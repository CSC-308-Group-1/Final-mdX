`timescale 1ns/1ps

`define SMEM_MAX 1024
`define RMEM_MAX 256
`define TRANSACTION_COUNT 5
`define DRIV_IF mem_intf.DriverInterface.Driver_cb
`define MON_IF mem_intf.ME_MONITOR.ME_monitor_cb
